module adder_tree_module
    #(
        parameter BITS  = 'd32,
        parameter CGES  = 'd49,
        parameter MAX   = $log2(CGES) + BITS,
        parameter INPUt = 'd7 
    )
    (
        input logic coeff
    );


    //adder block

endmodule